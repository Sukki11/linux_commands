module xor(a,b,c,res);
input a,b,c;
output res;
assign res=a^b;
endmodule


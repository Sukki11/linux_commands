module or(a,b,res);
input a,b;
output res;
assign res=a+b;
endmodule


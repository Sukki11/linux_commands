module



endmodule
